module foutbitbooth();
    
endmodule