module wallace_tb;
reg [31:0] a,b;
wire [63:0] product;

thirty_two_wallace_multipiler wallace(product[63:0],a[31:0],b[31:0]);

initial
begin
  $display("	WALLANCE MULTIPLIER (32 BIT)\n\n   ");
  $dumpfile("wallace_tb.vcd");
    // Module to capture and what level, 0 means all wires
    $dumpvars(0, wallace_tb);
end

initial
begin
      a=32'b00000000000000000000000000000000; b=32'b11111111111111111111111111111111;
  #30 a=32'b00000000000000000000000001111011; b=32'b00000000000000000000000101000001;
  #30 a=32'b00000000000000000000000100000000; b=32'b00000000000000000000000100000000;
  #30 a=32'b00000000011110000111100100110001; b=32'b00000000000000000000000000000010;
  #30 a=32'b00000000000000011000011010011111; b=32'b00000000000000000000111111111111; 
  #30 a=32'b11111111111111111111110101110010; b=32'b00000000000000000000000001111011; 
  #30 a=32'b00000000000000000000001010001110; b=32'b00000000000000000000000001111011; 
end

initial
begin
  $monitor(" %b * %b \n= %b \n\n (i.e %d * %d = %d) \n\n\n", a[31:0],b[31:0],product[63:0],a[31:0],b[31:0],product[63:0]); //(~a) + 1'b1
end


endmodule